package param_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    parameter PERIOD = 20;
    parameter SIZE   = 32;

endpackage :param_pkg