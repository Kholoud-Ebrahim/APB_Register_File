package rf_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    import seq_item_pkg::*;

    `include "rf_sequencer.svh"
    `include "rf_driver.svh"
    `include "rf_agent.svh"

endpackage :rf_agent_pkg