package seq_item_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    `include "rf_sequence_item.svh"

endpackage :seq_item_pkg