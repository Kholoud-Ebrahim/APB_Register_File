package test_lib_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    import rf_agent_pkg::*;
    import reg_model_pkg::*;
    import seq_lib_pkg::*;

    `include "apb_rf_env.svh"
        
    `include "apb_rf_base_test.svh"
    `include "rf_wr_ctl_test.svh"
    `include "rf_r_stat_test.svh"
    `include "rf_wr_to_test.svh"
    `include "rf_wr_t1_test.svh"

endpackage :test_lib_pkg