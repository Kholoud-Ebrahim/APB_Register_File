package apb_rf_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    import seq_item_pkg::*;
    
    import rf_agent_pkg::*;

    import reg_model_pkg::*;

    import seq_lib_pkg::*;


    import test_lib_pkg::*;
    
endpackage :apb_rf_pkg